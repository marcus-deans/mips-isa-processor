module or32(a,b,c);
  input [31:0]b;
  input [31:0]c;
  output [31:0]a;

  or o3233(a[0],b[0],c[0]);
  or o33244(a[1],b[1],c[1]);
  or o3325(a[2],b[2],c[2]);
  or o32263(a[3],b[3],c[3]);
  or o332973(a[4],b[4],c[4]);
  or o322338(a[5],b[5],c[5]);
  or o323398(a[6],b[6],c[6]);
  or o3383(a[7],b[7],c[7]);
  or o3322324(a[8],b[8],c[8]);
  or o33423(a[9],b[9],c[9]);
  or o3224323(a[10],b[10],c[10]);
  or o33723(a[11],b[11],c[11]);
  or o43323(a[12],b[12],c[12]);
  or o34323(a[13],b[13],c[13]);
  or o33653(a[14],b[14],c[14]);
  or o3772733(a[15],b[15],c[15]);
  or o366233(a[16],b[16],c[16]);
  or o3972933(a[17],b[17],c[17]);
  or o384323(a[18],b[18],c[18]);
  or o233323(a[19],b[19],c[19]);
  or o3422222333(a[20],b[20],c[20]);
  or o3324253(a[21],b[21],c[21]);
  or o34322233(a[22],b[22],c[22]);
  or o334553(a[23],b[23],c[23]);
  or o345323(a[24],b[24],c[24]);
  or o354226733(a[25],b[25],c[25]);
  or o33827653(a[26],b[26],c[26]);
  or o334253(a[27],b[27],c[27]);
  or o334563(a[28],b[28],c[28]);
  or o3334223(a[29],b[29],c[29]);
  or o334222663(a[30],b[30],c[30]);
  or o3223993(a[31],b[31],c[31]);
endmodule
