module and32(a,b,c);
  input [31:0]b;
  input [31:0]c;
  output [31:0]a;

  and o33t3(a[0],b[0],c[0]);
  and ot99(a[1],b[1],c[1]);
  and o33t5(a[2],b[2],c[2]);
  and o36t3(a[3],b[3],c[3]);
  and o33t73(a[4],b[4],c[4]);
  and o33t38(a[5],b[5],c[5]);
  and o333t98(a[6],b[6],c[6]);
  and o338tt3(a[7],b[7],c[7]);
  and o3t334(a[8],b[8],c[8]);
  and o334t3(a[9],b[9],c[9]);
  and o34t33(a[10],b[10],c[10]);
  and o336373(a[11],b[11],c[11]);
  and o43t33(a[12],b[12],c[12]);
  and o34876tr33(a[13],b[13],c[13]);
  and o33t653(a[14],b[14],c[14]);
  and o377733(a[15],b[15],c[15]);
  and o366t33(a[16],b[16],c[16]);
  and o397t933(a[17],b[17],c[17]);
  and o384t33(a[18],b[18],c[18]);
  and o233t33(a[19],b[19],c[19]);
  and o3433t3(a[20],b[20],c[20]);
  and o3345t3(a[21],b[21],c[21]);
  and o34t333(a[22],b[22],c[22]);
  and o33t4553(a[23],b[23],c[23]);
  and o345t33(a[24],b[24],c[24]);
  and o354t6733(a[25],b[25],c[25]);
  and o338t7653(a[26],b[26],c[26]);
  and o334t53(a[27],b[27],c[27]);
  and o334t563(a[28],b[28],c[28]);
  and o333t43(a[29],b[29],c[29]);
  and o334t663(a[30],b[30],c[30]);
  and o33t993(a[31],b[31],c[31]);
endmodule
