module bit32_not(out, a);
    input [31:0] a;
    output [31:0] out;

    not bit0(out[0], a[0]);
    not bit1(out[1], a[1]);
    not bit2(out[2], a[2]);
    not bit3(out[3], a[3]);
    not bit4(out[4], a[4]);
    not bit5(out[5], a[5]);
    not bit6(out[6], a[6]);
    not bit7(out[7], a[7]);
    not bit8(out[8], a[8]);
    not bit9(out[9], a[9]);
    not bit10(out[10], a[10]);
    not bit11(out[11], a[11]);
    not bit12(out[12], a[12]);
    not bit13(out[13], a[13]);
    not bit14(out[14], a[14]);
    not bit15(out[15], a[15]);
    not bit16(out[16], a[16]);
    not bit17(out[17], a[17]);
    not bit18(out[18], a[18]);
    not bit19(out[19], a[19]);
    not bit20(out[20], a[20]);
    not bit21(out[21], a[21]);
    not bit22(out[22], a[22]);
    not bit23(out[23], a[23]);
    not bit24(out[24], a[24]);
    not bit25(out[25], a[25]);
    not bit26(out[26], a[26]);
    not bit27(out[27], a[27]);
    not bit28(out[28], a[28]);
    not bit29(out[29], a[29]);
    not bit30(out[30], a[30]);
    not bit31(out[31], a[31]);

endmodule
