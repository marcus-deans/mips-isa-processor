module not32(a,b);
  input [31:0]b;
  output [31:0]a;

  not a3393(a[0],b[0]);
  not a339944(a[1],b[1]);
  not a3395(a[2],b[2]);
  not a3963(a[3],b[3]);
  not a399373(a[4],b[4]);
  not a93338(a[5],b[5]);
  not a933398(a[6],b[6]);
  not a93383(a[7],b[7]);
  not a33934(a[8],b[8]);
  not a33943(a[9],b[9]);
  not a3433(a[10],b[10]);
  not a3373(a[11],b[11]);
  not a4333(a[12],b[12]);
  not a34633(a[13],b[13]);
  not a33653(a[14],b[14]);
  not a377733(a[15],b[15]);
  not a36633(a[16],b[16]);
  not a397933(a[17],b[17]);
  not a38433(a[18],b[18]);
  not a23333(a[19],b[19]);
  not a34333(a[20],b[20]);
  not a55555(a[21],b[21]);
  not a3433553(a[22],b[22]);
  not a334553(a[23],b[23]);
  not a34533(a[24],b[24]);
  not a3546733(a[25],b[25]);
  not a3387653(a[26],b[26]);
  not a33453(a[27],b[27]);
  not a334563(a[28],b[28]);
  not a33343(a[29],b[29]);
  not a334663(a[30],b[30]);
  not a33993(a[31],b[31]);
endmodule
