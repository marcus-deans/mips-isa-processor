module decoder32(wr, enable, out);
    input [4:0] wr;
    input enable;

    output [31:0] out;

    // assign out = enable << wr;
    // wire [31:0] shifter_in;

    wire [31:0] validated;
    wire [4:0] n_wr;

    not NOT_0(n_wr[0], wr[0]);
    not NOT_1(n_wr[1], wr[1]);
    not NOT_2(n_wr[2], wr[2]);
    not NOT_3(n_wr[3], wr[3]);
    not NOT_4(n_wr[4], wr[4]);

    and decode0_gate(out[0], n_wr[4], n_wr[3], n_wr[2], n_wr[1], n_wr[0]);
    and decode1_gate(out[1], n_wr[4], n_wr[3], n_wr[2], n_wr[1], wr[0]);

    and decode2_gate(out[2], n_wr[4], n_wr[3], n_wr[2], wr[1], n_wr[0]);
    and decode3_gate(out[3], n_wr[4], n_wr[3], n_wr[2], wr[1], wr[0]);

    and decode4_gate(out[4], n_wr[4], n_wr[3], wr[2], n_wr[1], n_wr[0]);
    and decode5_gate(out[5], n_wr[4], n_wr[3], wr[2], n_wr[1], wr[0]);
    and decode6_gate(out[6], n_wr[4], n_wr[3], wr[2], wr[1], n_wr[0]);
    and decode7_gate(out[7], n_wr[4], n_wr[3], wr[2], wr[1], wr[0]);

    and decode8_gate(out[8], n_wr[4], wr[3], n_wr[2], n_wr[1], n_wr[0]);
    and decode9_gate(out[9], n_wr[4], wr[3], n_wr[2], n_wr[1], wr[0]);
    and decode10_gate(out[10], n_wr[4], wr[3], n_wr[2], wr[1], n_wr[0]);
    and decode11_gate(out[11], n_wr[4], wr[3], n_wr[2], wr[1], wr[0]);
    and decode12_gate(out[12], n_wr[4], wr[3], wr[2], n_wr[1], n_wr[0]);
    and decode13_gate(out[13], n_wr[4], wr[3], wr[2], n_wr[1], wr[0]);
    and decode14_gate(out[14], n_wr[4], wr[3], wr[2], wr[1], n_wr[0]);
    and decode15_gate(out[15], n_wr[4], wr[3], wr[2], wr[1], wr[0]);
    
    and decode16_gate(out[16], wr[4], n_wr[3], n_wr[2], n_wr[1], n_wr[0]);
    and decode17_gate(out[17], wr[4], n_wr[3], n_wr[2], n_wr[1], wr[0]);

    and decode18_gate(out[18], wr[4], n_wr[3], n_wr[2], wr[1], n_wr[0]);
    and decode19_gate(out[19], wr[4], n_wr[3], n_wr[2], wr[1], wr[0]);

    and decode20_gate(out[20], wr[4], n_wr[3], wr[2], n_wr[1], n_wr[0]);
    and decode21_gate(out[21], wr[4], n_wr[3], wr[2], n_wr[1], wr[0]);
    and decode22_gate(out[22], wr[4], n_wr[3], wr[2], wr[1], n_wr[0]);
    and decode23_gate(out[23], wr[4], n_wr[3], wr[2], wr[1], wr[0]);
    
    and decode24_gate(out[24], wr[4], wr[3], n_wr[2], n_wr[1], n_wr[0]);
    and decode25_gate(out[25], wr[4], wr[3], n_wr[2], n_wr[1], wr[0]);
    and decode26_gate(out[26], wr[4], wr[3], n_wr[2], wr[1], n_wr[0]);
    and decode27_gate(out[27], wr[4], wr[3], n_wr[2], wr[1], wr[0]);
    and decode28_gate(out[28], wr[4], wr[3], wr[2], n_wr[1], n_wr[0]);
    and decode29_gate(out[29], wr[4], wr[3], wr[2], n_wr[1], wr[0]);
    and decode30_gate(out[30], wr[4], wr[3], wr[2], wr[1], n_wr[0]);
    and decode31_gate(out[31], wr[4], wr[3], wr[2], wr[1], wr[0]);

    // and validate1_gate(validated[0], wr, 5'b00000);
    // and validate2_gate(validated[1], wr, 5'b00001);
    // and validate3_gate(validated[2], wr, 5'b00010);
    // and validate4_gate(validated[3], wr, 5'b00011);
    // and validate5_gate(validated[4], wr, 5'b00100);
    // and validate6_gate(validated[5], wr, 5'b00101);
    // and validate7_gate(validated[6], wr, 5'b00110);
    // and validate8_gate(validated[7], wr, 5'b00111);
    // and validate9_gate(validated[8], wr, 5'b01000);
    // and validate10_gate(validated[9], wr, 5'b01001);
    // and validate11_gate(validated[10], wr, 5'b01010);
    // and validate12_gate(validated[11], wr, 5'b01011);
    // and validate13_gate(validated[12], wr, 5'b01100);
    // and validate14_gate(validated[13], wr, 5'b01101);
    // and validate15_gate(validated[14], wr, 5'b01110);
    // and validate16_gate(validated[15], wr, 5'b01111);
    // and validate17_gate(validated[16], wr, 5'b10000);
    // and validate18_gate(validated[17], wr, 5'b10001);
    // and validate19_gate(validated[18], wr, 5'b10010);
    // and validate20_gate(validated[19], wr, 5'b10011);
    // and validate21_gate(validated[20], wr, 5'b10100);
    // and validate22_gate(validated[21], wr, 5'b10101);
    // and validate23_gate(validated[22], wr, 5'b10110);
    // and validate24_gate(validated[23], wr, 5'b10111);
    // and validate25_gate(validated[24], wr, 5'b11000);
    // and validate26_gate(validated[25], wr, 5'b11001);
    // and validate27_gate(validated[26], wr, 5'b11010);
    // and validate28_gate(validated[27], wr, 5'b11011);
    // and validate29_gate(validated[28], wr, 5'b11100);
    // and validate30_gate(validated[29], wr, 5'b11101);
    // and validate31_gate(validated[30], wr, 5'b11110);
    // and validate32_gate(validated[31], wr, 5'b11111);

    // and writeEnable0_gate(writeEnable[0], decoded[0], ctrl_writeEnable);
	// and writeEnable1_gate(writeEnable[1], decoded[1], ctrl_writeEnable);
	// and writeEnable2_gate(writeEnable[2], decoded[2], ctrl_writeEnable);
	// and writeEnable3_gate(writeEnable[3], decoded[3], ctrl_writeEnable);
	// and writeEnable4_gate(writeEnable[4], decoded[4], ctrl_writeEnable);
	// and writeEnable5_gate(writeEnable[5], decoded[5], ctrl_writeEnable);
	// and writeEnable6_gate(writeEnable[6], decoded[6], ctrl_writeEnable);
	// and writeEnable7_gate(writeEnable[7], decoded[7], ctrl_writeEnable);
	// and writeEnable8_gate(writeEnable[8], decoded[8], ctrl_writeEnable);
	// and writeEnable9_gate(writeEnable[9], decoded[9], ctrl_writeEnable);
	// and writeEnable10_gate(writeEnable[10], decoded[10], ctrl_writeEnable);
	// and writeEnable11_gate(writeEnable[11], decoded[11], ctrl_writeEnable);
	// and writeEnable12_gate(writeEnable[12], decoded[12], ctrl_writeEnable);
	// and writeEnable13_gate(writeEnable[13], decoded[13], ctrl_writeEnable);
	// and writeEnable14_gate(writeEnable[14], decoded[14], ctrl_writeEnable);
	// and writeEnable15_gate(writeEnable[15], decoded[15], ctrl_writeEnable);
	// and writeEnable16_gate(writeEnable[16], decoded[16], ctrl_writeEnable);
	// and writeEnable17_gate(writeEnable[17], decoded[17], ctrl_writeEnable);
	// and writeEnable18_gate(writeEnable[18], decoded[18], ctrl_writeEnable);
	// and writeEnable19_gate(writeEnable[19], decoded[19], ctrl_writeEnable);
	// and writeEnable20_gate(writeEnable[20], decoded[20], ctrl_writeEnable);
	// and writeEnable21_gate(writeEnable[21], decoded[21], ctrl_writeEnable);
	// and writeEnable22_gate(writeEnable[22], decoded[22], ctrl_writeEnable);
	// and writeEnable23_gate(writeEnable[23], decoded[23], ctrl_writeEnable);
	// and writeEnable24_gate(writeEnable[24], decoded[24], ctrl_writeEnable);
	// and writeEnable25_gate(writeEnable[25], decoded[25], ctrl_writeEnable);
	// and writeEnable26_gate(writeEnable[26], decoded[26], ctrl_writeEnable);
	// and writeEnable27_gate(writeEnable[27], decoded[27], ctrl_writeEnable);
	// and writeEnable28_gate(writeEnable[28], decoded[28], ctrl_writeEnable);
	// and writeEnable29_gate(writeEnable[29], decoded[29], ctrl_writeEnable);
	// and writeEnable30_gate(writeEnable[30], decoded[30], ctrl_writeEnable);
	// and writeEnable31_gate(writeEnable[31], decoded[31], ctrl_writeEnable);

    // assign out[0] = enable ? validated[0] : 1'b0;
    // assign out[1] = enable ? validated[1] : 1'b0;
    // assign out[2] = enable ? validated[2] : 1'b0;
    // assign out[3] = enable ? validated[3] : 1'b0;
    // assign out[4] = enable ? validated[4] : 1'b0;
    // assign out[5] = enable ? validated[5] : 1'b0;
    // assign out[6] = enable ? validated[6] : 1'b0;
    // assign out[7] = enable ? validated[7] : 1'b0;
    // assign out[8] = enable ? validated[8] : 1'b0;
    // assign out[9] = enable ? validated[9] : 1'b0;
    // assign out[10] = enable ? validated[10] : 1'b0;
    // assign out[11] = enable ? validated[11] : 1'b0;
    // assign out[12] = enable ? validated[12] : 1'b0;
    // assign out[13] = enable ? validated[13] : 1'b0;
    // assign out[14] = enable ? validated[14] : 1'b0;
    // assign out[15] = enable ? validated[15] : 1'b0;
    // assign out[16] = enable ? validated[16] : 1'b0;
    // assign out[17] = enable ? validated[17] : 1'b0;
    // assign out[18] = enable ? validated[18] : 1'b0;
    // assign out[19] = enable ? validated[19] : 1'b0;
    // assign out[20] = enable ? validated[20] : 1'b0;
    // assign out[21] = enable ? validated[21] : 1'b0;
    // assign out[22] = enable ? validated[22] : 1'b0;
    // assign out[23] = enable ? validated[23] : 1'b0;
    // assign out[24] = enable ? validated[24] : 1'b0;
    // assign out[25] = enable ? validated[25] : 1'b0;
    // assign out[26] = enable ? validated[26] : 1'b0;
    // assign out[27] = enable ? validated[27] : 1'b0;
    // assign out[28] = enable ? validated[28] : 1'b0;
    // assign out[29] = enable ? validated[29] : 1'b0;
    // assign out[30] = enable ? validated[30] : 1'b0;
    // assign out[31] = enable ? validated[31] : 1'b0;

    // and out0_gate(out[0], validated[0], enable);
    // and out1_gate(out[1], validated[1], enable);
    // and out2_gate(out[2], validated[2], enable);
    // and out3_gate(out[3], validated[3], enable);
    // and out4_gate(out[4], validated[4], enable);
    // and out5_gate(out[5], validated[5], enable);
    // and out6_gate(out[6], validated[6], enable);
    // and out7_gate(out[7], validated[7], enable);
    // and out8_gate(out[8], validated[8], enable);
    // and out9_gate(out[9], validated[9], enable);
    // and out10_gate(out[10], validated[10], enable);
    // and out11_gate(out[11], validated[11], enable);
    // and out12_gate(out[12], validated[12], enable);
    // and out13_gate(out[13], validated[13], enable);
    // and out14_gate(out[14], validated[14], enable);
    // and out15_gate(out[15], validated[15], enable);
    // and out16_gate(out[16], validated[16], enable);
    // and out17_gate(out[17], validated[17], enable);
    // and out18_gate(out[18], validated[18], enable);
    // and out19_gate(out[19], validated[19], enable);
    // and out20_gate(out[20], validated[20], enable);
    // and out21_gate(out[21], validated[21], enable);
    // and out22_gate(out[22], validated[22], enable);
    // and out23_gate(out[23], validated[23], enable);
    // and out24_gate(out[24], validated[24], enable);
    // and out25_gate(out[25], validated[25], enable);
    // and out26_gate(out[26], validated[26], enable);
    // and out27_gate(out[27], validated[27], enable);
    // and out28_gate(out[28], validated[28], enable);
    // and out29_gate(out[29], validated[29], enable);
    // and out30_gate(out[30], validated[30], enable);
    // and out31_gate(out[31], validated[31], enable);
endmodule